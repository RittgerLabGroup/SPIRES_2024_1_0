netcdf mod09ga_061_spi_h08v05_20240101.v2024.1.0 {
dimensions:
	time = UNLIMITED ; // (1 currently)
	x = 2400 ;
	y = 2400 ;
variables:
	double time(time) ;
		time:standard_name = "time" ;
		time:calendar = "standard" ;
		time:coverage_content_type = "coordinate" ;
		time:long_name = "ANSI date" ;
		time:units = "days since 2000-01-01 00:00:00" ;
		time:axis = "T" ;
		time:valid_range = 0., 1.79769313486232e+308 ;
    time:_Storage = "chunked" ;
		time:_ChunkSizes = 512 ;
		time:_Endianness = "little" ;
	double x(x) ;
		x:standard_name = "projection_x_coordinate" ;
		x:coverage_content_type = "coordinate" ;
		x:long_name = "x" ;
		x:units = "meters" ;
		x:axis = "X" ;
		x:valid_range = -20015109.3557974, 20015109.3557974 ;
    x:_Storage = "contiguous" ;
		x:_Endianness = "little" ;
	double y(y) ;
		y:standard_name = "projection_y_coordinate" ;
		y:coverage_content_type = "coordinate" ;
		y:long_name = "y" ;
		y:units = "meters" ;
		y:axis = "Y" ;
		y:valid_range = -10007554.6778987, 10007554.6778987 ;
    x:_Storage = "contiguous" ;
		x:_Endianness = "little" ;
	ubyte viewable_snow_fraction(time, y, x) ;
		viewable_snow_fraction:snowtoday_id = 54. ;
		viewable_snow_fraction:snowtoday_name = "viewable_snow_fraction_s" ;
		viewable_snow_fraction:long_name = "SPIReS-MODIS Terra viewable snow fraction" ;
		viewable_snow_fraction:units = "%" ;
		viewable_snow_fraction:_FillValue = 255UB ;
		viewable_snow_fraction:valid_range = 0UB, 100UB ;
		viewable_snow_fraction:comment = "Snow fraction from surface reflectance visible from satellite. Expressed in percent for each pixel, fillValue 255." ;
		viewable_snow_fraction:grid_mapping = "crs" ;
		viewable_snow_fraction:standard_name = "snow_area_fraction_viewable_from_above" ;
    viewable_snow_fraction:_Storage = "chunked" ;
		viewable_snow_fraction:_ChunkSizes = 1, 2400, 2400 ;
		viewable_snow_fraction:_DeflateLevel = 1 ;
		viewable_snow_fraction:_Shuffle = "true" ;
	ushort grain_size(time, y, x) ;
		grain_size:snowtoday_id = 57. ;
		grain_size:snowtoday_name = "grain_size_s" ;
		grain_size:long_name = "SPIReS-MODIS Terra grain size" ;
		grain_size:units = "um" ;
		grain_size:_FillValue = 65535US ;
		grain_size:valid_range = 40US, 1190US ;
		grain_size:comment = "Optical snow grain size based on SPIReS spectral mixture analysis. Expressed in micrometers for each pixel, fillValue 65535." ;
		grain_size:grid_mapping = "crs" ;
		grain_size:standard_name = "snow_grain_size" ;
    grain_size:_Storage = "chunked" ;
		grain_size:_ChunkSizes = 1, 2400, 2400 ;
		grain_size:_DeflateLevel = 1 ;
		grain_size:_Shuffle = "true" ;
	ushort dust_concentration(time, y, x) ;
		dust_concentration:snowtoday_id = 58. ;
		dust_concentration:snowtoday_name = "dust_concentration_s" ;
		dust_concentration:long_name = "SPIReS-MODIS Terra dust concentration" ;
		dust_concentration:units = "dppm" ;
		dust_concentration:_FillValue = 65535US ;
		dust_concentration:valid_range = 0US, 9500US ;
		dust_concentration:comment = "Dust concentration based on Spires spectral mixture analysis. Expressed in 10-7 unitless (or tenths of ppm) for each pixel, fillValue 65535." ;
		dust_concentration:grid_mapping = "crs" ;
    dust_concentration:_Storage = "chunked" ;
		dust_concentration:_ChunkSizes = 1, 2400, 2400 ;
		dust_concentration:_DeflateLevel = 1 ;
		dust_concentration:_Shuffle = "true" ;
	ubyte snow_fraction(time, y, x) ;
		snow_fraction:snowtoday_id = 55. ;
		snow_fraction:snowtoday_name = "snow_fraction_s" ;
		snow_fraction:long_name = "SPIReS-MODIS Terra on the ground snow fraction" ;
		snow_fraction:units = "%" ;
		snow_fraction:_FillValue = 255UB ;
		snow_fraction:valid_range = 0UB, 100UB ;
		snow_fraction:comment = "Viewable snow fraction adjusted using a Geometrical Optical model. Expressed in percent of pixel, for each pixel, fillValue 255." ;
		snow_fraction:grid_mapping = "crs" ;
		snow_fraction:standard_name = "surface_snow_area_fraction" ;
    snow_fraction:_Storage = "chunked" ;
		snow_fraction:_ChunkSizes = 1, 2400, 2400 ;
		snow_fraction:_DeflateLevel = 1 ;
		snow_fraction:_Shuffle = "true" ;
	ushort snow_cover_duration(time, y, x) ;
		snow_cover_duration:snowtoday_id = 61. ;
		snow_cover_duration:snowtoday_name = "snow_cover_days_s" ;
		snow_cover_duration:long_name = "SPIReS-MODIS Terra snow cover duration" ;
		snow_cover_duration:units = "day" ;
		snow_cover_duration:_FillValue = 65535US ;
		snow_cover_duration:valid_range = 0US, 366US ;
		snow_cover_duration:comment = "The number of days since the start of the water year with a value greater than the threshold for viewable snow cover fraction, for each pixel. Water year N is set from 10/1/(N – 1) to 9/30/N for the northern hemisphere, and from 4/1/(N – 1) to 3/31/N for the southern hemisphere. Expressed in days for each pixel, fillValue 65535." ;
		snow_cover_duration:grid_mapping = "crs" ;
    snow_cover_duration:_Storage = "chunked" ;
		snow_cover_duration:_ChunkSizes = 1, 2400, 2400 ;
		snow_cover_duration:_DeflateLevel = 1 ;
		snow_cover_duration:_Shuffle = "true" ;
	ubyte albedo(time, y, x) ;
		albedo:snowtoday_id = 62. ;
		albedo:snowtoday_name = "albedo_s" ;
		albedo:long_name = "SPIReS-MODIS Terra snow albedo assuming flat surface darkened by light-absorbing particles" ;
		albedo:units = "%" ;
		albedo:_FillValue = 255UB ;
		albedo:valid_range = 0UB, 100UB ;
		albedo:comment = "Spires reflected fraction of broadband (0.28-4.00 micrometer) solar radiation, based on optical grain size accounting for darkening by light-absorbing impurities, no adjustment to account for slope and aspect of the terrain. Expressed in percent for each pixel, fillValue 255." ;
		albedo:grid_mapping = "crs" ;
    albedo:_Storage = "chunked" ;
		albedo:_ChunkSizes = 1, 2400, 2400 ;
		albedo:_DeflateLevel = 1 ;
		albedo:_Shuffle = "true" ;
	ushort radiative_forcing(time, y, x) ;
		radiative_forcing:snowtoday_id = 63. ;
		radiative_forcing:snowtoday_name = "radiative_forcing_s" ;
		radiative_forcing:long_name = "SPIReS-MODIS Terra radiative forcing on snow" ;
		radiative_forcing:units = "W m-2" ;
		radiative_forcing:_FillValue = 65535US ;
		radiative_forcing:valid_range = 0US, 500US ;
		radiative_forcing:comment = "Additional energy absorbed by the snowpack from light-absorbing impurities assuming a clear sky. Expressed in Watt per square meter for each pixel, fillValue 65535." ;
		radiative_forcing:grid_mapping = "crs" ;
		radiative_forcing:standard_name = "surface_downward_heat_flux_in_snow" ;
    radiative_forcing:_Storage = "chunked" ;
		radiative_forcing:_ChunkSizes = 1, 2400, 2400 ;
		radiative_forcing:_DeflateLevel = 1 ;
		radiative_forcing:_Shuffle = "true" ;
	ubyte deltavis(time, y, x) ;
		deltavis:snowtoday_id = 96. ;
		deltavis:snowtoday_name = "deltavis_s" ;
		deltavis:long_name = "SPIReS-MODIS Terra decrease in snow albedo from light absorbing particles" ;
		deltavis:units = "%" ;
		deltavis:_FillValue = 255UB ;
		deltavis:valid_range = 0UB, 75UB ;
		deltavis:comment = "Decrease in observed visible broadband (0.350-0.876 micrometer) albedo estimated using SPIReS-MODIS Terra retrieved snow grain size and dust concentration. Expressed in percent for each pixel, fillValue 255." ;
		deltavis:grid_mapping = "crs" ;
    deltavis:_Storage = "chunked" ;
		deltavis:_ChunkSizes = 1, 2400, 2400 ;
		deltavis:_DeflateLevel = 1 ;
		deltavis:_Shuffle = "true" ;
	ubyte albedo_muZ(time, y, x) ;
		albedo_muZ:snowtoday_id = 99. ;
		albedo_muZ:snowtoday_name = "albedo_muZ_s" ;
		albedo_muZ:long_name = "SPIReS-MODIS Terra snow albedo on slope darkened by light-absorbing particles, typically dust." ;
		albedo_muZ:units = "%" ;
		albedo_muZ:_FillValue = 255UB ;
		albedo_muZ:valid_range = 0UB, 100UB ;
		albedo_muZ:comment = "Spires reflected fraction of broadband (0.28-4.00 micrometer) solar radiation, based on optical grain size accounting for darkening by light-absorbing impurities, adjusted to account for slope and aspect of the terrain. Expressed in percent for each pixel, fillValue 255." ;
		albedo_muZ:grid_mapping = "crs" ;
    albedo_muZ:_Storage = "chunked" ;
		albedo_muZ:_ChunkSizes = 1, 2400, 2400 ;
		albedo_muZ:_DeflateLevel = 1 ;
		albedo_muZ:_Shuffle = "true" ;
	char crs ;
		crs:grid_mapping_name = "sinusoidal" ;
		crs:false_easting = 0. ;
		crs:false_northing = 0. ;
		crs:longitude_of_projection_origin = 0. ;
		crs:longitude_of_central_meridian = 0. ;
		crs:long_name = "Sinusoidal projection definition" ;
		crs:longitude_of_prime_meridian = 0. ;
		crs:semi_major_axis = 6371007.181 ;
		crs:inverse_flattening = 0. ;
		crs:proj4 = "+proj=sinu +lon_0=0 +x_0=0 +y_0=0 +a=6371007.181 +b=6371007.181 +units=m +no_defs +nadgrids=@null +wktext" ;
		crs:spatial_ref = "PROJCS[\"MODIS Sinusoidal\",GEOGCS[\"User with datum World Geodetic Survey 1984\",DATUM[\"unnamed\",SPHEROID[\"unnamed\",6371007.181,0]],PRIMEM[\"Greenwich\",0],UNIT[\"degree\",0.0174532925199433,AUTHORITY[\"EPSG\",\"9122\"]]],PROJECTION[\"Sinusoidal\"],PARAMETER[\"longitude_of_center\",0],PARAMETER[\"false_easting\",0],PARAMETER[\"false_northing\",0],UNIT[\"metre\",1,AUTHORITY[\"EPSG\",\"9001\"]],AXIS[\"Easting\",EAST],AXIS[\"Northing\",NORTH]]" ;
		crs:crs_wkt = "PROJCS[\"MODIS Sinusoidal\",GEOGCS[\"User with datum World Geodetic Survey 1984\",DATUM[\"unnamed\",SPHEROID[\"unnamed\",6371007.181,0]],PRIMEM[\"Greenwich\",0],UNIT[\"degree\",0.0174532925199433,AUTHORITY[\"EPSG\",\"9122\"]]],PROJECTION[\"Sinusoidal\"],PARAMETER[\"longitude_of_center\",0],PARAMETER[\"false_easting\",0],PARAMETER[\"false_northing\",0],UNIT[\"metre\",1,AUTHORITY[\"EPSG\",\"9001\"]],AXIS[\"Easting\",EAST],AXIS[\"Northing\",NORTH]]" ;
		crs:GeoTransform = "-11119505.19766523316502571106 463.31271656938469050147 0.0 4447802.07906609307974576950 0.0 -463.31271656938469050147 " ;
    crs:_Storage = "contiguous" ;

// global attributes:
    :id = "TO BE UPDATED" ;
		:title = "MODIS/Terra L3 Daily 500m SIN Grid SPIReS Snow Cover, Snow Albedo, and other Snow Physical Properties, Version v2024.hist." ;
    :citation = "Mandatory citation for any work, including articles, reports, presentations, abstracts and posters as: Rittger, K., S. J. P. Lenard, R. T. Palomaki, E. H. Bair, and J. Dozier. 2024. MODIS/Terra L3 Daily 500m SIN Grid SPIReS Snow Cover, Snow Albedo, and other Snow Physical Properties, Version v2024.1.0. INSTAAR, University of Colorado, Boulder, CO, USA. Digital Media. [@TO UPDATE DOI THERE]. https://github.com/sebastien-lenard/snow-today.   https://nsidc.org/snow-today." ;
    :license = "Creative Commons BY 4.0. You are free to (1) share: copy and redistribute the material in any medium or format for any purpose, even commercially; (2) Adapt: remix, transform, and build upon the material for any purpose, even commercially; Under the following terms, (3) Attribution: You must give appropriate credit, provide a link to the license, and indicate if changes were made. You may do so in any reasonable manner, but not in any way that suggests the licensor endorses you or your use. https://creativecommons.org/licenses/by/4.0/." ;
		:summary = "This dataset contains daily raster images of snow cover and snow surface properties. Snow cover, grain size and dust concentration were unmixed from the daily reflectance of the MOD09GA Terra Collection 6 v061 (Vermote and Wolfe, 2021) using an adapted version of the SPIReS algorithm (Bair et al., 2021), that we named SPIReS v2024.1.0, with a removal of clouds and data errors. The data were then temporally interpolated to fill the cloudy days, and the snow cover duration was calculated from the start of the water year (October 1st for the northern hemisphere, April 1st for the southern one). Deltavis, radiative forcing, and albedos were calculated using an adaptation of the ParBal algorithm (Bair et al., 2018), that we included in SPIReS v2024.hist." ;
		:source = "MOD09GA Terra Collection 6 v061" ;
		:comment = "Snow cover validated with 3 m airborne snow maps on 116 days (Stillinger et al., 2023); Snow albedo validated using terrain correct in-situ observations at 3 sites for ~20 years with spatial comparisons to 31 ASO Inc hyperspectral airborne flights (Palomaki et al., RSE, in review). Preliminary radiative forcing evaluation performed at 1 site in the San Juan mountains of Colorado." ;
		:metadata_link = "TO BE UPDATED" ;
		:product_version = "v2024.1.0" ;
		:software_version_id = "c196e7d" ;
		:publisher_institution = "Institute for Arctic and Alpine Research" ;
		:publisher_name = "Institute for Arctic and Alpine Research" ;
		:publisher_type = "institution" ;
		:publisher_url = "https://nsidc.org/snow-today" ;
		:publisher_email = "snow-today@nsidc.org" ;
		:Conventions = "CF-1.10, ACDD-1.3" ;
		:standard_name_vocabulary = "CF Standard Name Table (v82, 06 July 2023)" ;
		:history = "" ;
		:references = "Bair, E.H., T. Stillinger, and J. Dozier. 2021. Snow Property Inversion from Remote Sensing (SPIReS): A generalized multispectral unmixing approach with examples from MODIS and Landsat 8 OLI. IEEE Transactions on Geoscience and Remote Sensing 59.9: 7270-7284, doi: 10.1109/TGRS.2020.3040328. https://github.com/edwardbair/SPIRES. Palomaki, R., K. Rittger, S.J.P, Lenard, E.H, Bair, J., Dozier, M. Skiles, and T.H. Painter (in revision). Assessment for mapping snow albedo from MODIS. Remote Sensing of Environment. Stillinger, T., K. Rittger, M.S. Raleigh, A. Michell, R.E. Davis, and E.H. Bair. 2023. Landsat, MODIS, and VIIRS snow cover mapping algorithm performance as validated by airborne lidar datasets. The Cryosphere 17: 567-590, doi: 10.5194/tc-17-567-2023. Bair, E. H., A. Abreu Calfa, K. Rittger, and J. Dozier. 2018. Using machine learning for real-time estimates of snow water equivalent in the watersheds of Afghanistan. The Cryosphere 12.5: 1579-1594, doi: 10.5194/tc-12-1579-2018. https://github.com/edwardbair/ParBal. Bair, E. H., K. Rittger, R. E. Davis, T. H. Painter, and Dozier, J. 2016. Validating reconstruction of snow water equivalent in California\'s Sierra Nevada using measurements from the NASA Airborne Snow Observatory. Water Resources Research 52, doi: 10.1002/2016WR018704. Rittger, K., Bair, E.H., Kahl, A., and Dozier, J. 2016. Spatial estimates of snow water equivalent from reconstruction. Advances in Water Resources 94: 345-363, doi: 10.1016/j.advwatres.2016.05.015. Vermote, E., and R. Wolfe. 2021. MODIS/Terra Surface Reflectance Daily L2G Global 1km and 500m SIN Grid V061. Distributed by NASA EOSDIS Land Processes Distributed Active Archive Center, doi: 10.5067/MODIS/MOD09GA.061.MODIS." ;
		:acknowledgement = "These data are produced and supported by the Institute of Arctic and Alpine Research. The data products were produced with funding from NASA grants 80NSSC22K0703 (Rittger, TAS), 80NSSC20K1721 (Rittger, HMA), 80NSSC22K0929 (Rittger, WR), 80NSSC23K1456 (Rittger, Alps), 80NSSC24K1270 (Rittger, IDS). This work utilized the Alpine high performance computing resource at the University of Colorado Boulder. Alpine is jointly funded by the University of Colorado Boulder, the University of Colorado Anschutz, and Colorado State University. Data storage supported by the University of Colorado Boulder PetaLibrary." ;
		:creator_name = "Karl Rittger" ;
		:creator_url = "https://www.colorado.edu/instaar/karl-rittger" ;
		:creator_email = "karl.rittger@colorado.edu" ;
		:contributor_name = "Karl Rittger, Sebastien J. P. Lenard, Ross T. Palomaki" ;
		:contributor_role = "principal_investigator, research_scientist, research_scientist" ;
		:geospatial_bounds_crs = "EPSG:4326" ;
		:geospatial_bounds = "POLYGON((40.00000000 -130.54072893, 40.00000000 -117.48665604, 30.00000000 -103.92304845, 30.00000000 -115.47005384, 40.00000000 -130.54072893))" ;
		:time_coverage_start = "2024-01-01T00:00:00.000+0000" ;
		:time_coverage_end = "2024-01-02T00:00:00.000+0000" ;
		:time_coverage_duration = "P0Y0M1DT0H0M0S" ;
    :versionOf_SPIReS = "v2024.1.0" ;
    :versionOf_SPIReS_alternative = "v2024.0d" ;
		:date_created = "2024-12-06T23:54:48+00:00" ;
		:date_modified = "2024-12-06T23:54:48+00:00" ;
    :_NCProperties = "version=2,netcdf=4.7.4,hdf5=1.8.12" ;
		:_SuperblockVersion = 0 ;
		:_IsNetcdf4 = 1 ;
		:_Format = "netCDF-4" ;
}
